module glfw3

pub enum GLFWKey {
    key_a = C.GLFW_KEY_A
    key_b = C.GLFW_KEY_B
    key_c = C.GLFW_KEY_C
    key_d = C.GLFW_KEY_D
    key_e = C.GLFW_KEY_E
    key_f = C.GLFW_KEY_F
    key_g = C.GLFW_KEY_G
    key_h = C.GLFW_KEY_H
    key_i = C.GLFW_KEY_I
    key_j = C.GLFW_KEY_J
    key_k = C.GLFW_KEY_K
    key_l = C.GLFW_KEY_L
    key_m = C.GLFW_KEY_M
    key_n = C.GLFW_KEY_N
    key_o = C.GLFW_KEY_O
    key_p = C.GLFW_KEY_P
    key_q = C.GLFW_KEY_Q
    key_r = C.GLFW_KEY_R
    key_s = C.GLFW_KEY_S
    key_t = C.GLFW_KEY_T
    key_u = C.GLFW_KEY_U
    key_v = C.GLFW_KEY_V
    key_w = C.GLFW_KEY_W
    key_x = C.GLFW_KEY_X
    key_y = C.GLFW_KEY_Y
    key_z = C.GLFW_KEY_Z
    key_0 = C.GLFW_KEY_0
    key_1 = C.GLFW_KEY_1
    key_2 = C.GLFW_KEY_2
    key_3 = C.GLFW_KEY_3
    key_4 = C.GLFW_KEY_4
    key_5 = C.GLFW_KEY_5
    key_6 = C.GLFW_KEY_6
    key_7 = C.GLFW_KEY_7
    key_8 = C.GLFW_KEY_8
    key_9 = C.GLFW_KEY_9
    key_f1 = C.GLFW_KEY_F1
    key_f2 = C.GLFW_KEY_F2
    key_f3 = C.GLFW_KEY_F3
    key_f4 = C.GLFW_KEY_F4
    key_f5 = C.GLFW_KEY_F5
    key_f6 = C.GLFW_KEY_F6
    key_f7 = C.GLFW_KEY_F7
    key_f8 = C.GLFW_KEY_F8
    key_f9 = C.GLFW_KEY_F9
    key_f10 = C.GLFW_KEY_F10
    key_f11 = C.GLFW_KEY_F11
    key_f12 = C.GLFW_KEY_F12
    key_right = C.GLFW_KEY_RIGHT
    key_left = C.GLFW_KEY_LEFT
    key_down = C.GLFW_KEY_DOWN
    key_up = C.GLFW_KEY_UP
    key_apostrophe = C.GLFW_KEY_APOSTROPHE
    key_backslash = C.GLFW_KEY_BACKSLASH
    key_backspace = C.GLFW_KEY_BACKSPACE
    key_caps_lock = C.GLFW_KEY_CAPS_LOCK
    key_comma = C.GLFW_KEY_COMMA
    key_delete = C.GLFW_KEY_DELETE
    key_end = C.GLFW_KEY_END
    key_enter = C.GLFW_KEY_ENTER
    key_equal = C.GLFW_KEY_EQUAL
    key_escape = C.GLFW_KEY_ESCAPE
    key_grave_accent = C.GLFW_KEY_GRAVE_ACCENT
    key_home = C.GLFW_KEY_HOME
    key_insert = C.GLFW_KEY_INSERT
    key_last = C.GLFW_KEY_LAST
    key_left_alt = C.GLFW_KEY_LEFT_ALT
    key_left_bracket = C.GLFW_KEY_LEFT_BRACKET
    key_left_control = C.GLFW_KEY_LEFT_CONTROL
    key_left_shift = C.GLFW_KEY_LEFT_SHIFT
    key_left_super = C.GLFW_KEY_LEFT_SUPER
    key_menu = C.GLFW_KEY_MENU
    key_minus = C.GLFW_KEY_MINUS
    key_num_lock = C.GLFW_KEY_NUM_LOCK
    key_page_down = C.GLFW_KEY_PAGE_DOWN
    key_page_up = C.GLFW_KEY_PAGE_UP
    key_period = C.GLFW_KEY_PERIOD
    key_right_alt = C.GLFW_KEY_RIGHT_ALT
    key_right_bracket = C.GLFW_KEY_RIGHT_BRACKET
    key_right_control = C.GLFW_KEY_RIGHT_CONTROL
    key_right_shift = C.GLFW_KEY_RIGHT_SHIFT
    key_right_super = C.GLFW_KEY_RIGHT_SUPER
    key_scroll_lock = C.GLFW_KEY_SCROLL_LOCK
    key_semicolon = C.GLFW_KEY_SEMICOLON
    key_slash = C.GLFW_KEY_SLASH
    key_space = C.GLFW_KEY_SPACE
    key_tab = C.GLFW_KEY_TAB
    key_kp_add = C.GLFW_KEY_KP_ADD
    key_kp_decimal = C.GLFW_KEY_KP_DECIMAL
    key_kp_divide = C.GLFW_KEY_KP_DIVIDE
    key_kp_enter = C.GLFW_KEY_KP_ENTER
    key_kp_equal = C.GLFW_KEY_KP_EQUAL
    key_kp_multiply = C.GLFW_KEY_KP_MULTIPLY
    key_kp_subtract = C.GLFW_KEY_KP_SUBTRACT
    key_kp_0 = C.GLFW_KEY_KP_0
    key_kp_1 = C.GLFW_KEY_KP_1
    key_kp_2 = C.GLFW_KEY_KP_2
    key_kp_3 = C.GLFW_KEY_KP_3
    key_kp_4 = C.GLFW_KEY_KP_4
    key_kp_5 = C.GLFW_KEY_KP_5
    key_kp_6 = C.GLFW_KEY_KP_6
    key_kp_7 = C.GLFW_KEY_KP_7
    key_kp_8 = C.GLFW_KEY_KP_8
    key_kp_9 = C.GLFW_KEY_KP_9
}
