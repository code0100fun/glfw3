module glfw3

#flag -DGLFW_INCLUDE_NONE
#flag -lglfw3

#include <GLFW/glfw3.h>
