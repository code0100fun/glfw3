module glfw3

#flag -DGLFW_INCLUDE_NONE
#flag windows -lglfw3
#flag linux -lglfw

#include <GLFW/glfw3.h>
